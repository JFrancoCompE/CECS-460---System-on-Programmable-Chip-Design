`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/15/2020 08:30:27 PM
// Design Name: 
// Module Name: ADRS_DECODE
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ADRS_DECODE(
    input write_strobe,
    input read_strobe,
    input port_id_15,
    input [2:0] port_id,
    output [7:0] read,
    output [7:0] write
    );
    
    //always@(*)
      //  if(port_id_15 && write_strobe)
    
    
endmodule
